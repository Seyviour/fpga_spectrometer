module i2s_clk_gen (
    input wire clk_in,
    output wire i2s_clk
);
    //VENDOR SPECIFIC
endmodule